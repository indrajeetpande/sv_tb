class or_mon;

endclass
