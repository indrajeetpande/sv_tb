class or_sco;
endclass
