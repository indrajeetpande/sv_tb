`include "and_gate.v"
`include "base_pkt.sv"
`include "interface.sv"
`include "generator.sv"
`include "driver.sv"
`include "mon.sv"
`include "sco.sv"
`include "env.sv"
`include "test.sv"
`include "top.sv"
