interface and_inf;
    bit a;
    bit b;
    bit y;
endinterface
